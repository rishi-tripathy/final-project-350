/******************************************************************************
 *                                                                            *
 * Module:       Hexadecimal_To_Seven_Segment                                 *
 * Description:                                                               *
 *      This module converts hexadecimal numbers for seven segment displays.  *
 *                                                                            *
 ******************************************************************************/

module Decimal_To_Seven_Segment (
	// Inputs
	clk,
	dec_number,

	// Bidirectional

	// Outputs
	seven_seg_display_ones,
	seven_seg_display_tens
);

/*****************************************************************************
 *                           Parameter Declarations                          *
 *****************************************************************************/


/*****************************************************************************
 *                             Port Declarations                             *
 *****************************************************************************/
// Inputs
input clk;
input		[7:0]	dec_number;

reg[3:0] ones, tens;

always @(posedge clk) begin

	ones <= dec_number % 4'd10;
	tens <= dec_number / 4'd10;
end

 

// Bidirectional

// Outputs
output		[6:0]	seven_seg_display_ones;
output		[6:0]	seven_seg_display_tens;


/*****************************************************************************
 *                            Combinational Logic                            *
 *****************************************************************************/

assign seven_seg_display_ones =
		({7{(ones == 4'h0)}} & 7'b1000000) |
		({7{(ones == 4'h1)}} & 7'b1111001) |
		({7{(ones == 4'h2)}} & 7'b0100100) |
		({7{(ones == 4'h3)}} & 7'b0110000) |
		({7{(ones == 4'h4)}} & 7'b0011001) |
		({7{(ones == 4'h5)}} & 7'b0010010) |
		({7{(ones == 4'h6)}} & 7'b0000010) |
		({7{(ones == 4'h7)}} & 7'b1111000) |
		({7{(ones == 4'h8)}} & 7'b0000000) |
		({7{(ones == 4'h9)}} & 7'b0010000) |
		({7{(ones == 4'hA)}} & 7'b0001000) |
		({7{(ones == 4'hB)}} & 7'b0000011) |
		({7{(ones == 4'hC)}} & 7'b1000110) |
		({7{(ones == 4'hD)}} & 7'b0100001) |
		({7{(ones == 4'hE)}} & 7'b0000110) |
		({7{(ones == 4'hF)}} & 7'b0001110); 

		
assign seven_seg_display_tens =
		({7{(tens == 4'h0)}} & 7'b1000000) |
		({7{(tens == 4'h1)}} & 7'b1111001) |
		({7{(tens == 4'h2)}} & 7'b0100100) |
		({7{(tens == 4'h3)}} & 7'b0110000) |
		({7{(tens == 4'h4)}} & 7'b0011001) |
		({7{(tens == 4'h5)}} & 7'b0010010) |
		({7{(tens == 4'h6)}} & 7'b0000010) |
		({7{(tens == 4'h7)}} & 7'b1111000) |
		({7{(tens == 4'h8)}} & 7'b0000000) |
		({7{(tens == 4'h9)}} & 7'b0010000) |
		({7{(tens == 4'hA)}} & 7'b0001000) |
		({7{(tens == 4'hB)}} & 7'b0000011) |
		({7{(tens == 4'hC)}} & 7'b1000110) |
		({7{(tens == 4'hD)}} & 7'b0100001) |
		({7{(tens == 4'hE)}} & 7'b0000110) |
		({7{(tens == 4'hF)}} & 7'b0001110); 


/*****************************************************************************
 *                              Internal Modules                             *
 *****************************************************************************/


endmodule

