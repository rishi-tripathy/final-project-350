module mw_pipeline(ir, result, q_dmem, out, data_mw, ir_q, clk, en, clr, exception, exception_q);

	input [31:0] ir, result, q_dmem;
	output [31:0] data_mw, ir_q, out;
	input clk, en, clr, exception;
	output exception_q;
	
	dffe_ref dff00(.d(exception), .q(exception_q), .clr(clr), .clk(clk), .en(en));
	
	dffe_ref dff0a(.d(q_dmem[0]), .q(data_mw[0]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1a(.d(q_dmem[1]), .q(data_mw[1]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2a(.d(q_dmem[2]), .q(data_mw[2]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff3a(.d(q_dmem[3]), .q(data_mw[3]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff4a(.d(q_dmem[4]), .q(data_mw[4]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff5a(.d(q_dmem[5]), .q(data_mw[5]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff6a(.d(q_dmem[6]), .q(data_mw[6]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff7a(.d(q_dmem[7]), .q(data_mw[7]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff8a(.d(q_dmem[8]), .q(data_mw[8]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff9a(.d(q_dmem[9]), .q(data_mw[9]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1a0(.d(q_dmem[10]), .q(data_mw[10]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1a1(.d(q_dmem[11]), .q(data_mw[11]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1a2(.d(q_dmem[12]), .q(data_mw[12]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1a3(.d(q_dmem[13]), .q(data_mw[13]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1a4(.d(q_dmem[14]), .q(data_mw[14]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1a5(.d(q_dmem[15]), .q(data_mw[15]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1a6(.d(q_dmem[16]), .q(data_mw[16]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1a7(.d(q_dmem[17]), .q(data_mw[17]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1a8(.d(q_dmem[18]), .q(data_mw[18]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1a9(.d(q_dmem[19]), .q(data_mw[19]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2a0(.d(q_dmem[20]), .q(data_mw[20]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2a1(.d(q_dmem[21]), .q(data_mw[21]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2a2(.d(q_dmem[22]), .q(data_mw[22]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2a3(.d(q_dmem[23]), .q(data_mw[23]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2a4(.d(q_dmem[24]), .q(data_mw[24]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2a5(.d(q_dmem[25]), .q(data_mw[25]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2a6(.d(q_dmem[26]), .q(data_mw[26]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2a7(.d(q_dmem[27]), .q(data_mw[27]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2a8(.d(q_dmem[28]), .q(data_mw[28]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2a9(.d(q_dmem[29]), .q(data_mw[29]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff3a0(.d(q_dmem[30]), .q(data_mw[30]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff3a1(.d(q_dmem[31]), .q(data_mw[31]), .clr(clr), .clk(clk), .en(en));

	dffe_ref dff0(.d(result[0]), .q(out[0]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1(.d(result[1]), .q(out[1]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2(.d(result[2]), .q(out[2]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff3(.d(result[3]), .q(out[3]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff4(.d(result[4]), .q(out[4]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff5(.d(result[5]), .q(out[5]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff6(.d(result[6]), .q(out[6]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff7(.d(result[7]), .q(out[7]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff8(.d(result[8]), .q(out[8]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff9(.d(result[9]), .q(out[9]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff10(.d(result[10]), .q(out[10]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff11(.d(result[11]), .q(out[11]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff12(.d(result[12]), .q(out[12]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff13(.d(result[13]), .q(out[13]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff14(.d(result[14]), .q(out[14]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff15(.d(result[15]), .q(out[15]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff16(.d(result[16]), .q(out[16]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff17(.d(result[17]), .q(out[17]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff18(.d(result[18]), .q(out[18]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff19(.d(result[19]), .q(out[19]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff20(.d(result[20]), .q(out[20]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff21(.d(result[21]), .q(out[21]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff22(.d(result[22]), .q(out[22]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff23(.d(result[23]), .q(out[23]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff24(.d(result[24]), .q(out[24]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff25(.d(result[25]), .q(out[25]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff26(.d(result[26]), .q(out[26]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff27(.d(result[27]), .q(out[27]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff28(.d(result[28]), .q(out[28]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff29(.d(result[29]), .q(out[29]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff30(.d(result[30]), .q(out[30]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff31(.d(result[31]), .q(out[31]), .clr(clr), .clk(clk), .en(en));
	
	dffe_ref dff0b(.d(ir[0]), .q(ir_q[0]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1b(.d(ir[1]), .q(ir_q[1]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2b(.d(ir[2]), .q(ir_q[2]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff3b(.d(ir[3]), .q(ir_q[3]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff4b(.d(ir[4]), .q(ir_q[4]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff5b(.d(ir[5]), .q(ir_q[5]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff6b(.d(ir[6]), .q(ir_q[6]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff7b(.d(ir[7]), .q(ir_q[7]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff8b(.d(ir[8]), .q(ir_q[8]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff9b(.d(ir[9]), .q(ir_q[9]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1b0(.d(ir[10]), .q(ir_q[10]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1b1(.d(ir[11]), .q(ir_q[11]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1b2(.d(ir[12]), .q(ir_q[12]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1b3(.d(ir[13]), .q(ir_q[13]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1b4(.d(ir[14]), .q(ir_q[14]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1b5(.d(ir[15]), .q(ir_q[15]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1b6(.d(ir[16]), .q(ir_q[16]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1b7(.d(ir[17]), .q(ir_q[17]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1b8(.d(ir[18]), .q(ir_q[18]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff1b9(.d(ir[19]), .q(ir_q[19]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2b0(.d(ir[20]), .q(ir_q[20]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2b1(.d(ir[21]), .q(ir_q[21]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2b2(.d(ir[22]), .q(ir_q[22]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2b3(.d(ir[23]), .q(ir_q[23]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2b4(.d(ir[24]), .q(ir_q[24]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2b5(.d(ir[25]), .q(ir_q[25]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2b6(.d(ir[26]), .q(ir_q[26]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2b7(.d(ir[27]), .q(ir_q[27]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2b8(.d(ir[28]), .q(ir_q[28]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff2b9(.d(ir[29]), .q(ir_q[29]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff3b0(.d(ir[30]), .q(ir_q[30]), .clr(clr), .clk(clk), .en(en));
	dffe_ref dff3b1(.d(ir[31]), .q(ir_q[31]), .clr(clr), .clk(clk), .en(en));

endmodule
